module top_module (
    output out);
     assign out = 1'b00;
endmodule
